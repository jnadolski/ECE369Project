`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// ECE369A - Computer Architecture
// Laboratory  1
// Module - InstructionMemory.v
// Description - 32-Bit wide instruction memory.
//
// INPUT:-
// Address: 32-Bit address input port.
//
// OUTPUT:-
// Instruction: 32-Bit output port.
//
// FUNCTIONALITY:-
// Similar to the DataMemory, this module should also be byte-addressed
// (i.e., ignore bits 0 and 1 of 'Address'). All of the instructions will be 
// hard-coded into the instruction memory, so there is no need to write to the 
// InstructionMemory.  The contents of the InstructionMemory is the machine 
// language program to be run on your MIPS processor.
//
//
//we will store the machine code for a code written in C later. for now initialize 
//each entry to be its index * 3 (memory[i] = i * 3;)
//all you need to do is give an address as input and read the contents of the 
//address on your output port. 
// 
//Using a 32bit address you will index into the memory, output the contents of that specific 
//address. for data memory we are using 1K word of storage space. for the instruction memory 
//you may assume smaller size for practical purpose. you can use 128 words as the size and 
//hardcode the values.  in this case you need 7 bits to index into the memory. 
//
//be careful with the least two significant bits of the 32bit address. those help us index 
//into one of the 4 bytes in a word. therefore you will need to use bit [8-2] of the input address. 


////////////////////////////////////////////////////////////////////////////////

module InstructionMemory(Address, Instruction); 

    input [31:0] Address;        // Input Address 

    output reg [31:0] Instruction;    // Instruction at memory location Address
    
    reg [31:0] memory [512:0];
    integer i;
    
    initial begin
//    for(i=0; i<127;i=i+1) begin
//    memory[i] = i*3;
//    end

//memory[0] <= 32'b00100000000100000000000000000001;
//memory[1] <= 32'b00000000000000000000000000000000;
//memory[2] <= 32'b00000000000000000000000000000000;
//memory[3] <= 32'b00000000000000000000000000000000;
//memory[4] <= 32'b00000000000000000000000000000000;
//memory[5] <= 32'b00000000000000000000000000000000;
//memory[6] <= 32'b00100000000100010000000000000001;
//memory[7] <= 32'b00000000000000000000000000000000;
//memory[8] <= 32'b00000000000000000000000000000000;
//memory[9] <= 32'b00000000000000000000000000000000;
//memory[10] <= 32'b00000000000000000000000000000000;
//memory[11] <= 32'b00000000000000000000000000000000;
//memory[12] <= 32'b00000010000100011000000000100100;
//memory[13] <= 32'b00000000000000000000000000000000;
//memory[14] <= 32'b00000000000000000000000000000000;
//memory[15] <= 32'b00000000000000000000000000000000;
//memory[16] <= 32'b00000000000000000000000000000000;
//memory[17] <= 32'b00000000000000000000000000000000;
//memory[18] <= 32'b00000010000000001000000000100100;
//memory[19] <= 32'b00000000000000000000000000000000;
//memory[20] <= 32'b00000000000000000000000000000000;
//memory[21] <= 32'b00000000000000000000000000000000;
//memory[22] <= 32'b00000000000000000000000000000000;
//memory[23] <= 32'b00000000000000000000000000000000;
//memory[24] <= 32'b00000010001100001000000000100010;
//memory[25] <= 32'b00000000000000000000000000000000;
//memory[26] <= 32'b00000000000000000000000000000000;
//memory[27] <= 32'b00000000000000000000000000000000;
//memory[28] <= 32'b00000000000000000000000000000000;
//memory[29] <= 32'b00000000000000000000000000000000;
//memory[30] <= 32'b00000010000000001000000000100111;
//memory[31] <= 32'b00000000000000000000000000000000;
//memory[32] <= 32'b00000000000000000000000000000000;
//memory[33] <= 32'b00000000000000000000000000000000;
//memory[34] <= 32'b00000000000000000000000000000000;
//memory[35] <= 32'b00000000000000000000000000000000;
//memory[36] <= 32'b00000010000000001000000000100111;
//memory[37] <= 32'b00000000000000000000000000000000;
//memory[38] <= 32'b00000000000000000000000000000000;
//memory[39] <= 32'b00000000000000000000000000000000;
//memory[40] <= 32'b00000000000000000000000000000000;
//memory[41] <= 32'b00000000000000000000000000000000;
//memory[42] <= 32'b00000000000000001000000000100101;
//memory[43] <= 32'b00000000000000000000000000000000;
//memory[44] <= 32'b00000000000000000000000000000000;
//memory[45] <= 32'b00000000000000000000000000000000;
//memory[46] <= 32'b00000000000000000000000000000000;
//memory[47] <= 32'b00000000000000000000000000000000;
//memory[48] <= 32'b00000010001000001000000000100101;
//memory[49] <= 32'b00000000000000000000000000000000;
//memory[50] <= 32'b00000000000000000000000000000000;
//memory[51] <= 32'b00000000000000000000000000000000;
//memory[52] <= 32'b00000000000000000000000000000000;
//memory[53] <= 32'b00000000000000000000000000000000;
//memory[54] <= 32'b00000000000100001000000010000000;
//memory[55] <= 32'b00000000000000000000000000000000;
//memory[56] <= 32'b00000000000000000000000000000000;
//memory[57] <= 32'b00000000000000000000000000000000;
//memory[58] <= 32'b00000000000000000000000000000000;
//memory[59] <= 32'b00000000000000000000000000000000;
//memory[60] <= 32'b00000010001100001000000000000100;
//memory[61] <= 32'b00000000000000000000000000000000;
//memory[62] <= 32'b00000000000000000000000000000000;
//memory[63] <= 32'b00000000000000000000000000000000;
//memory[64] <= 32'b00000000000000000000000000000000;
//memory[65] <= 32'b00000000000000000000000000000000;
//memory[66] <= 32'b00000010000000001000000000101010;
//memory[67] <= 32'b00000000000000000000000000000000;
//memory[68] <= 32'b00000000000000000000000000000000;
//memory[69] <= 32'b00000000000000000000000000000000;
//memory[70] <= 32'b00000000000000000000000000000000;
//memory[71] <= 32'b00000000000000000000000000000000;
//memory[72] <= 32'b00000010000100011000000000101010;
//memory[73] <= 32'b00000000000000000000000000000000;
//memory[74] <= 32'b00000000000000000000000000000000;
//memory[75] <= 32'b00000000000000000000000000000000;
//memory[76] <= 32'b00000000000000000000000000000000;
//memory[77] <= 32'b00000000000000000000000000000000;
//memory[78] <= 32'b00000000000100011000000001000011;
//memory[79] <= 32'b00000000000000000000000000000000;
//memory[80] <= 32'b00000000000000000000000000000000;
//memory[81] <= 32'b00000000000000000000000000000000;
//memory[82] <= 32'b00000000000000000000000000000000;
//memory[83] <= 32'b00000000000000000000000000000000;
//memory[84] <= 32'b00000000000100011000000000000111;
//memory[85] <= 32'b00000000000000000000000000000000;
//memory[86] <= 32'b00000000000000000000000000000000;
//memory[87] <= 32'b00000000000000000000000000000000;
//memory[88] <= 32'b00000000000000000000000000000000;
//memory[89] <= 32'b00000000000000000000000000000000;
//memory[90] <= 32'b00000000000100011000000001000010;
//memory[91] <= 32'b00000000000000000000000000000000;
//memory[92] <= 32'b00000000000000000000000000000000;
//memory[93] <= 32'b00000000000000000000000000000000;
//memory[94] <= 32'b00000000000000000000000000000000;
//memory[95] <= 32'b00000000000000000000000000000000;
//memory[96] <= 32'b00000000000100011000000011000000;
//memory[97] <= 32'b00000000000000000000000000000000;
//memory[98] <= 32'b00000000000000000000000000000000;
//memory[99] <= 32'b00000000000000000000000000000000;
//memory[100] <= 32'b00000000000000000000000000000000;
//memory[101] <= 32'b00000000000000000000000000000000;
//memory[102] <= 32'b00000000000100001000000011000010;
//memory[103] <= 32'b00000000000000000000000000000000;
//memory[104] <= 32'b00000000000000000000000000000000;
//memory[105] <= 32'b00000000000000000000000000000000;
//memory[106] <= 32'b00000000000000000000000000000000;
//memory[107] <= 32'b00000000000000000000000000000000;
//memory[108] <= 32'b00000010001100001000000000000100;
//memory[109] <= 32'b00000000000000000000000000000000;
//memory[110] <= 32'b00000000000000000000000000000000;
//memory[111] <= 32'b00000000000000000000000000000000;
//memory[112] <= 32'b00000000000000000000000000000000;
//memory[113] <= 32'b00000000000000000000000000000000;
//memory[114] <= 32'b00000010001100001000000000000110;
//memory[115] <= 32'b00000000000000000000000000000000;
//memory[116] <= 32'b00000000000000000000000000000000;
//memory[117] <= 32'b00000000000000000000000000000000;
//memory[118] <= 32'b00000000000000000000000000000000;
//memory[119] <= 32'b00000000000000000000000000000000;
//memory[120] <= 32'b00000010000100011000000000100110;
//memory[121] <= 32'b00000000000000000000000000000000;
//memory[122] <= 32'b00000000000000000000000000000000;
//memory[123] <= 32'b00000000000000000000000000000000;
//memory[124] <= 32'b00000000000000000000000000000000;
//memory[125] <= 32'b00000000000000000000000000000000;
//memory[126] <= 32'b00000010000100011000000000100110;
//memory[127] <= 32'b00000000000000000000000000000000;
//memory[128] <= 32'b00000000000000000000000000000000;
//memory[129] <= 32'b00000000000000000000000000000000;
//memory[130] <= 32'b00000000000000000000000000000000;
//memory[131] <= 32'b00000000000000000000000000000000;
//memory[132] <= 32'b00100000000100100000000000000100;
//memory[133] <= 32'b00000000000000000000000000000000;
//memory[134] <= 32'b00000000000000000000000000000000;
//memory[135] <= 32'b00000000000000000000000000000000;
//memory[136] <= 32'b00000000000000000000000000000000;
//memory[137] <= 32'b00000000000000000000000000000000;
//memory[138] <= 32'b01110010000100101000000000000010;
//memory[139] <= 32'b00000000000000000000000000000000;
//memory[140] <= 32'b00000000000000000000000000000000;
//memory[141] <= 32'b00000000000000000000000000000000;
//memory[142] <= 32'b00000000000000000000000000000000;
//memory[143] <= 32'b00000000000000000000000000000000;
//memory[144] <= 32'b00100010000100000000000000000100;
//memory[145] <= 32'b00000000000000000000000000000000;
//memory[146] <= 32'b00000000000000000000000000000000;
//memory[147] <= 32'b00000000000000000000000000000000;
//memory[148] <= 32'b00000000000000000000000000000000;
//memory[149] <= 32'b00000000000000000000000000000000;
//memory[150] <= 32'b00110010000100000000000000000000;
//memory[151] <= 32'b00000000000000000000000000000000;
//memory[152] <= 32'b00000000000000000000000000000000;
//memory[153] <= 32'b00000000000000000000000000000000;
//memory[154] <= 32'b00000000000000000000000000000000;
//memory[155] <= 32'b00000000000000000000000000000000;
//memory[156] <= 32'b00110110000100000000000000000001;
//memory[157] <= 32'b00000000000000000000000000000000;
//memory[158] <= 32'b00000000000000000000000000000000;
//memory[159] <= 32'b00000000000000000000000000000000;
//memory[160] <= 32'b00000000000000000000000000000000;
//memory[161] <= 32'b00000000000000000000000000000000;
//memory[162] <= 32'b00101010000100000000000000000000;
//memory[163] <= 32'b00000000000000000000000000000000;
//memory[164] <= 32'b00000000000000000000000000000000;
//memory[165] <= 32'b00000000000000000000000000000000;
//memory[166] <= 32'b00000000000000000000000000000000;
//memory[167] <= 32'b00000000000000000000000000000000;
//memory[168] <= 32'b00101010000100000000000000000001;
//memory[169] <= 32'b00000000000000000000000000000000;
//memory[170] <= 32'b00000000000000000000000000000000;
//memory[171] <= 32'b00000000000000000000000000000000;
//memory[172] <= 32'b00000000000000000000000000000000;
//memory[173] <= 32'b00000000000000000000000000000000;
//memory[174] <= 32'b00111010000100000000000000000001;
//memory[175] <= 32'b00000000000000000000000000000000;
//memory[176] <= 32'b00000000000000000000000000000000;
//memory[177] <= 32'b00000000000000000000000000000000;
//memory[178] <= 32'b00000000000000000000000000000000;
//memory[179] <= 32'b00000000000000000000000000000000;
//memory[180] <= 32'b00111010000100000000000000000001;
//memory[181] <= 32'b00000000000000000000000000000000;
//memory[182] <= 32'b00000000000000000000000000000000;
//memory[183] <= 32'b00000000000000000000000000000000;
//memory[184] <= 32'b00000000000000000000000000000000;
//memory[185] <= 32'b00000000000000000000000000000000;
//memory[186] <= 32'b00100000000100001111111111111110;
//memory[187] <= 32'b00000000000000000000000000000000;
//memory[188] <= 32'b00000000000000000000000000000000;
//memory[189] <= 32'b00000000000000000000000000000000;
//memory[190] <= 32'b00000000000000000000000000000000;
//memory[191] <= 32'b00000000000000000000000000000000;
//memory[192] <= 32'b00100000000100010000000000000010;
//memory[193] <= 32'b00000000000000000000000000000000;
//memory[194] <= 32'b00000000000000000000000000000000;
//memory[195] <= 32'b00000000000000000000000000000000;
//memory[196] <= 32'b00000000000000000000000000000000;
//memory[197] <= 32'b00000000000000000000000000000000;
//memory[198] <= 32'b00000010001100001001000000101011;
//memory[199] <= 32'b00000000000000000000000000000000;
//memory[200] <= 32'b00000000000000000000000000000000;
//memory[201] <= 32'b00000000000000000000000000000000;
//memory[202] <= 32'b00000000000000000000000000000000;
//memory[203] <= 32'b00000000000000000000000000000000;
//memory[204] <= 32'b00101110001100001111111111111110;
//memory[205] <= 32'b00000000000000000000000000000000;
//memory[206] <= 32'b00000000000000000000000000000000;
//memory[207] <= 32'b00000000000000000000000000000000;
//memory[208] <= 32'b00000000000000000000000000000000;
//memory[209] <= 32'b00000000000000000000000000000000;
//memory[210] <= 32'b00000010001000001000000000001010;
//memory[211] <= 32'b00000000000000000000000000000000;
//memory[212] <= 32'b00000000000000000000000000000000;
//memory[213] <= 32'b00000000000000000000000000000000;
//memory[214] <= 32'b00000000000000000000000000000000;
//memory[215] <= 32'b00000000000000000000000000000000;
//memory[216] <= 32'b00000000000100011000000000001011;
//memory[217] <= 32'b00000000000000000000000000000000;
//memory[218] <= 32'b00000000000000000000000000000000;
//memory[219] <= 32'b00000000000000000000000000000000;
//memory[220] <= 32'b00000000000000000000000000000000;
//memory[221] <= 32'b00000000000000000000000000000000;
//memory[222] <= 32'b00000010001100101000000000100000;
//memory[223] <= 32'b00000000000000000000000000000000;
//memory[224] <= 32'b00000000000000000000000000000000;
//memory[225] <= 32'b00000000000000000000000000000000;
//memory[226] <= 32'b00000000000000000000000000000000;
//memory[227] <= 32'b00000000000000000000000000000000;
//memory[228] <= 32'b00100000000100001111111111111110;
//memory[229] <= 32'b00000000000000000000000000000000;
//memory[230] <= 32'b00000000000000000000000000000000;
//memory[231] <= 32'b00000000000000000000000000000000;
//memory[232] <= 32'b00000000000000000000000000000000;
//memory[233] <= 32'b00000000000000000000000000000000;
//memory[234] <= 32'b00000010001100001000100000100001;
//memory[235] <= 32'b00000000000000000000000000000000;
//memory[236] <= 32'b00000000000000000000000000000000;
//memory[237] <= 32'b00000000000000000000000000000000;
//memory[238] <= 32'b00000000000000000000000000000000;
//memory[239] <= 32'b00000000000000000000000000000000;
//memory[240] <= 32'b00100100000100011111111111111111;
//memory[241] <= 32'b00000000000000000000000000000000;
//memory[242] <= 32'b00000000000000000000000000000000;
//memory[243] <= 32'b00000000000000000000000000000000;
//memory[244] <= 32'b00000000000000000000000000000000;
//memory[245] <= 32'b00000000000000000000000000000000;
//memory[246] <= 32'b00100000000100100000000000100000;
//memory[247] <= 32'b00000000000000000000000000000000;
//memory[248] <= 32'b00000000000000000000000000000000;
//memory[249] <= 32'b00000000000000000000000000000000;
//memory[250] <= 32'b00000000000000000000000000000000;
//memory[251] <= 32'b00000000000000000000000000000000;
//memory[252] <= 32'b00000010001100100000000000011000;
//memory[253] <= 32'b00000000000000000000000000000000;
//memory[254] <= 32'b00000000000000000000000000000000;
//memory[255] <= 32'b00000000000000000000000000000000;
//memory[256] <= 32'b00000000000000000000000000000000;
//memory[257] <= 32'b00000000000000000000000000000000;
//memory[258] <= 32'b00000000000000001010000000010000;
//memory[259] <= 32'b00000000000000000000000000000000;
//memory[260] <= 32'b00000000000000000000000000000000;
//memory[261] <= 32'b00000000000000000000000000000000;
//memory[262] <= 32'b00000000000000000000000000000000;
//memory[263] <= 32'b00000000000000000000000000000000;
//memory[264] <= 32'b00000000000000001010100000010010;
//memory[265] <= 32'b00000000000000000000000000000000;
//memory[266] <= 32'b00000000000000000000000000000000;
//memory[267] <= 32'b00000000000000000000000000000000;
//memory[268] <= 32'b00000000000000000000000000000000;
//memory[269] <= 32'b00000000000000000000000000000000;
//memory[270] <= 32'b00000010001100100000000000011001;
//memory[271] <= 32'b00000000000000000000000000000000;
//memory[272] <= 32'b00000000000000000000000000000000;
//memory[273] <= 32'b00000000000000000000000000000000;
//memory[274] <= 32'b00000000000000000000000000000000;
//memory[275] <= 32'b00000000000000000000000000000000;
//memory[276] <= 32'b00000000000000001010000000010000;
//memory[277] <= 32'b00000000000000000000000000000000;
//memory[278] <= 32'b00000000000000000000000000000000;
//memory[279] <= 32'b00000000000000000000000000000000;
//memory[280] <= 32'b00000000000000000000000000000000;
//memory[281] <= 32'b00000000000000000000000000000000;
//memory[282] <= 32'b00000000000000001010100000010010;
//memory[283] <= 32'b00000000000000000000000000000000;
//memory[284] <= 32'b00000000000000000000000000000000;
//memory[285] <= 32'b00000000000000000000000000000000;
//memory[286] <= 32'b00000000000000000000000000000000;
//memory[287] <= 32'b00000000000000000000000000000000;
//memory[288] <= 32'b01110010001100100000000000000000;
//memory[289] <= 32'b00000000000000000000000000000000;
//memory[290] <= 32'b00000000000000000000000000000000;
//memory[291] <= 32'b00000000000000000000000000000000;
//memory[292] <= 32'b00000000000000000000000000000000;
//memory[293] <= 32'b00000000000000000000000000000000;
//memory[294] <= 32'b00000000000000001010000000010000;
//memory[295] <= 32'b00000000000000000000000000000000;
//memory[296] <= 32'b00000000000000000000000000000000;
//memory[297] <= 32'b00000000000000000000000000000000;
//memory[298] <= 32'b00000000000000000000000000000000;
//memory[299] <= 32'b00000000000000000000000000000000;
//memory[300] <= 32'b00000000000000001010100000010010;
//memory[301] <= 32'b00000000000000000000000000000000;
//memory[302] <= 32'b00000000000000000000000000000000;
//memory[303] <= 32'b00000000000000000000000000000000;
//memory[304] <= 32'b00000000000000000000000000000000;
//memory[305] <= 32'b00000000000000000000000000000000;
//memory[306] <= 32'b00000010010000000000000000010001;
//memory[307] <= 32'b00000000000000000000000000000000;
//memory[308] <= 32'b00000000000000000000000000000000;
//memory[309] <= 32'b00000000000000000000000000000000;
//memory[310] <= 32'b00000000000000000000000000000000;
//memory[311] <= 32'b00000000000000000000000000000000;
//memory[312] <= 32'b00000010001000000000000000010011;
//memory[313] <= 32'b00000000000000000000000000000000;
//memory[314] <= 32'b00000000000000000000000000000000;
//memory[315] <= 32'b00000000000000000000000000000000;
//memory[316] <= 32'b00000000000000000000000000000000;
//memory[317] <= 32'b00000000000000000000000000000000;
//memory[318] <= 32'b00000000000000001010000000010000;
//memory[319] <= 32'b00000000000000000000000000000000;
//memory[320] <= 32'b00000000000000000000000000000000;
//memory[321] <= 32'b00000000000000000000000000000000;
//memory[322] <= 32'b00000000000000000000000000000000;
//memory[323] <= 32'b00000000000000000000000000000000;
//memory[324] <= 32'b00000000000000001010100000010010;
//memory[325] <= 32'b00000000000000000000000000000000;
//memory[326] <= 32'b00000000000000000000000000000000;
//memory[327] <= 32'b00000000000000000000000000000000;
//memory[328] <= 32'b00000000000000000000000000000000;
//memory[329] <= 32'b00000000000000000000000000000000;
//memory[330] <= 32'b00110010001100011111111111111111;
//memory[331] <= 32'b00000000000000000000000000000000;
//memory[332] <= 32'b00000000000000000000000000000000;
//memory[333] <= 32'b00000000000000000000000000000000;
//memory[334] <= 32'b00000000000000000000000000000000;
//memory[335] <= 32'b00000000000000000000000000000000;
//memory[336] <= 32'b01110010100100100000000000000100;
//memory[337] <= 32'b00000000000000000000000000000000;
//memory[338] <= 32'b00000000000000000000000000000000;
//memory[339] <= 32'b00000000000000000000000000000000;
//memory[340] <= 32'b00000000000000000000000000000000;
//memory[341] <= 32'b00000000000000000000000000000000;
//memory[342] <= 32'b00000000000000001010000000010000;
//memory[343] <= 32'b00000000000000000000000000000000;
//memory[344] <= 32'b00000000000000000000000000000000;
//memory[345] <= 32'b00000000000000000000000000000000;
//memory[346] <= 32'b00000000000000000000000000000000;
//memory[347] <= 32'b00000000000000000000000000000000;
//memory[348] <= 32'b00000000000000001010100000010010;
//memory[349] <= 32'b00000000000000000000000000000000;
//memory[350] <= 32'b00000000000000000000000000000000;
//memory[351] <= 32'b00000000000000000000000000000000;
//memory[352] <= 32'b00000000000000000000000000000000;
//memory[353] <= 32'b00000000000000000000000000000000;
//memory[354] <= 32'b00100000000100100000000000000001;
//memory[355] <= 32'b00000000000000000000000000000000;
//memory[356] <= 32'b00000000000000000000000000000000;
//memory[357] <= 32'b00000000000000000000000000000000;
//memory[358] <= 32'b00000000000000000000000000000000;
//memory[359] <= 32'b00000000000000000000000000000000;
//memory[360] <= 32'b00000000001100101000111111000010;
//memory[361] <= 32'b00000000000000000000000000000000;
//memory[362] <= 32'b00000000000000000000000000000000;
//memory[363] <= 32'b00000000000000000000000000000000;
//memory[364] <= 32'b00000000000000000000000000000000;
//memory[365] <= 32'b00000000000000000000000000000000;
//memory[366] <= 32'b00100000000101000000000000011111;
//memory[367] <= 32'b00000000000000000000000000000000;
//memory[368] <= 32'b00000000000000000000000000000000;
//memory[369] <= 32'b00000000000000000000000000000000;
//memory[370] <= 32'b00000000000000000000000000000000;
//memory[371] <= 32'b00000000000000000000000000000000;
//memory[372] <= 32'b00000010100100011000100001000110;
//memory[373] <= 32'b00000000000000000000000000000000;
//memory[374] <= 32'b00000000000000000000000000000000;
//memory[375] <= 32'b00000000000000000000000000000000;
//memory[376] <= 32'b00000000000000000000000000000000;
//memory[377] <= 32'b00000000000000000000000000000000;
//memory[378] <= 32'b00110100000100010000111111110000;
//memory[379] <= 32'b00000000000000000000000000000000;
//memory[380] <= 32'b00000000000000000000000000000000;
//memory[381] <= 32'b00000000000000000000000000000000;
//memory[382] <= 32'b00000000000000000000000000000000;
//memory[383] <= 32'b00000000000000000000000000000000;
//memory[384] <= 32'b01111100000100011010010000100000;
//memory[385] <= 32'b00000000000000000000000000000000;
//memory[386] <= 32'b00000000000000000000000000000000;
//memory[387] <= 32'b00000000000000000000000000000000;
//memory[388] <= 32'b00000000000000000000000000000000;
//memory[389] <= 32'b00000000000000000000000000000000;
//memory[390] <= 32'b01111100000100011010011000100000;
//memory[391] <= 32'b00000000000000000000000000000000;
//memory[392] <= 32'b00000000000000000000000000000000;
//memory[393] <= 32'b00000000000000000000000000000000;
//memory[394] <= 32'b00000000000000000000000000000000;
//memory[395] <= 32'b00000000000000000000000000000000;



// //LOAD/STORE TESTING AND BYTE ADDRESSING 
//memory[0] <= 32'b00111100000010001010101111001110;	//		lui	$t0, 43982
// memory[1] <= 32'b00000000000000000000000000000000;    //        nop
// memory[2] <= 32'b00000000000000000000000000000000;    //        nop
// memory[3] <= 32'b00000000000000000000000000000000;    //        nop
// memory[4] <= 32'b00000000000000000000000000000000;    //        nop
// memory[5] <= 32'b00000000000000000000000000000000;    //        nop
// memory[6] <= 32'b00100001000010001101110010111010;    //        addi    $t0, $t0, 56506
// memory[7] <= 32'b00000000000000000000000000000000;    //        nop
// memory[8] <= 32'b00000000000000000000000000000000;    //        nop
// memory[9] <= 32'b00000000000000000000000000000000;    //        nop
// memory[10] <= 32'b00000000000000000000000000000000;    //        nop
// memory[11] <= 32'b00000000000000000000000000000000;    //        nop
// memory[12] <= 32'b00100000000010010000000000000100;    //        addi    $t1, $0, 4
// memory[13] <= 32'b00000000000000000000000000000000;    //        nop
// memory[14] <= 32'b00000000000000000000000000000000;    //        nop
// memory[15] <= 32'b00000000000000000000000000000000;    //        nop
// memory[16] <= 32'b00000000000000000000000000000000;    //        nop
// memory[17] <= 32'b00000000000000000000000000000000;    //        nop
// memory[18] <= 32'b10101101001010000000000000000000;    //        sw    $t0, 0($t1)
// memory[19] <= 32'b00000000000000000000000000000000;    //        nop
// memory[20] <= 32'b00000000000000000000000000000000;    //        nop
// memory[21] <= 32'b00000000000000000000000000000000;    //        nop
// memory[22] <= 32'b00000000000000000000000000000000;    //        nop
// memory[23] <= 32'b00000000000000000000000000000000;    //        nop
// memory[24] <= 32'b10101101001010000000000000000100;    //        sw    $t0, 4($t1)
// memory[25] <= 32'b00000000000000000000000000000000;    //        nop
// memory[26] <= 32'b00000000000000000000000000000000;    //        nop
// memory[27] <= 32'b00000000000000000000000000000000;    //        nop
// memory[28] <= 32'b00000000000000000000000000000000;    //        nop
// memory[29] <= 32'b00000000000000000000000000000000;    //        nop
// memory[30] <= 32'b00100001001010010000000000001000;    //        addi    $t1, $t1, 8
// memory[31] <= 32'b00000000000000000000000000000000;    //        nop
// memory[32] <= 32'b00000000000000000000000000000000;    //        nop
// memory[33] <= 32'b00000000000000000000000000000000;    //        nop
// memory[34] <= 32'b00000000000000000000000000000000;    //        nop
// memory[35] <= 32'b00000000000000000000000000000000;    //        nop
// memory[36] <= 32'b10100101001010000000000000000000;    //        sh    $t0, 0($t1)
// memory[37] <= 32'b00000000000000000000000000000000;    //        nop
// memory[38] <= 32'b00000000000000000000000000000000;    //        nop
// memory[39] <= 32'b00000000000000000000000000000000;    //        nop
// memory[40] <= 32'b00000000000000000000000000000000;    //        nop
// memory[41] <= 32'b00000000000000000000000000000000;    //        nop
// memory[42] <= 32'b10100101001010000000000000000010;    //        sh    $t0, 2($t1)
// memory[43] <= 32'b00000000000000000000000000000000;    //        nop
// memory[44] <= 32'b00000000000000000000000000000000;    //        nop
// memory[45] <= 32'b00000000000000000000000000000000;    //        nop
// memory[46] <= 32'b00000000000000000000000000000000;    //        nop
// memory[47] <= 32'b00000000000000000000000000000000;    //        nop
// memory[48] <= 32'b00100001001010010000000000000100;    //        addi    $t1, $t1, 4
// memory[49] <= 32'b00000000000000000000000000000000;    //        nop
// memory[50] <= 32'b00000000000000000000000000000000;    //        nop
// memory[51] <= 32'b00000000000000000000000000000000;    //        nop
// memory[52] <= 32'b00000000000000000000000000000000;    //        nop
// memory[53] <= 32'b00000000000000000000000000000000;    //        nop
// memory[54] <= 32'b10100001001010000000000000000000;    //        sb    $t0, 0($t1)
// memory[55] <= 32'b00000000000000000000000000000000;    //        nop
// memory[56] <= 32'b00000000000000000000000000000000;    //        nop
// memory[57] <= 32'b00000000000000000000000000000000;    //        nop
// memory[58] <= 32'b00000000000000000000000000000000;    //        nop
// memory[59] <= 32'b00000000000000000000000000000000;    //        nop
// memory[60] <= 32'b10100001001010000000000000000010;    //        sb    $t0, 2($t1)
// memory[61] <= 32'b00000000000000000000000000000000;    //        nop
// memory[62] <= 32'b00000000000000000000000000000000;    //        nop
// memory[63] <= 32'b00000000000000000000000000000000;    //        nop
// memory[64] <= 32'b00000000000000000000000000000000;    //        nop
// memory[65] <= 32'b00000000000000000000000000000000;    //        nop
// memory[66] <= 32'b00100000000010010000000000000100;    //        addi    $t1, $0, 4
// memory[67] <= 32'b00000000000000000000000000000000;    //        nop
// memory[68] <= 32'b00000000000000000000000000000000;    //        nop
// memory[69] <= 32'b00000000000000000000000000000000;    //        nop
// memory[70] <= 32'b00000000000000000000000000000000;    //        nop
// memory[71] <= 32'b00000000000000000000000000000000;    //        nop
// memory[72] <= 32'b10001101001010100000000000000000;    //        lw    $t2, 0($t1)
// memory[73] <= 32'b00000000000000000000000000000000;    //        nop
// memory[74] <= 32'b00000000000000000000000000000000;    //        nop
// memory[75] <= 32'b00000000000000000000000000000000;    //        nop
// memory[76] <= 32'b00000000000000000000000000000000;    //        nop
// memory[77] <= 32'b00000000000000000000000000000000;    //        nop
// memory[78] <= 32'b10001101001010110000000000000100;    //        lw    $t3, 4($t1)
// memory[79] <= 32'b00000000000000000000000000000000;    //        nop
// memory[80] <= 32'b00000000000000000000000000000000;    //        nop
// memory[81] <= 32'b00000000000000000000000000000000;    //        nop
// memory[82] <= 32'b00000000000000000000000000000000;    //        nop
// memory[83] <= 32'b00000000000000000000000000000000;    //        nop
// memory[84] <= 32'b10000101001011000000000000000000;    //        lh    $t4, 0($t1)
// memory[85] <= 32'b00000000000000000000000000000000;    //        nop
// memory[86] <= 32'b00000000000000000000000000000000;    //        nop
// memory[87] <= 32'b00000000000000000000000000000000;    //        nop
// memory[88] <= 32'b00000000000000000000000000000000;    //        nop
// memory[89] <= 32'b00000000000000000000000000000000;    //        nop
// memory[90] <= 32'b10000101001011010000000000000010;    //        lh    $t5, 2($t1)
// memory[91] <= 32'b00000000000000000000000000000000;    //        nop
// memory[92] <= 32'b00000000000000000000000000000000;    //        nop
// memory[93] <= 32'b00000000000000000000000000000000;    //        nop
// memory[94] <= 32'b00000000000000000000000000000000;    //        nop
// memory[95] <= 32'b00000000000000000000000000000000;    //        nop
// memory[96] <= 32'b10000001001011100000000000000000;    //        lb    $t6, 0($t1)
// memory[97] <= 32'b00000000000000000000000000000000;    //        nop
// memory[98] <= 32'b00000000000000000000000000000000;    //        nop
// memory[99] <= 32'b00000000000000000000000000000000;    //        nop
// memory[100] <= 32'b00000000000000000000000000000000;    //        nop
// memory[101] <= 32'b00000000000000000000000000000000;    //        nop
// memory[102] <= 32'b10000001001011110000000000000010;    //        lb    $t7, 2($t1)


/* //JUMP TESTING 
memory[0] <= 32'b00100000000010000000000000001010;	//		addi	$t0, $0, 10
memory[1] <= 32'b00000000000000000000000000000000;	//		nop
memory[2] <= 32'b00000000000000000000000000000000;	//		nop
memory[3] <= 32'b00000000000000000000000000000000;	//		nop
memory[4] <= 32'b00000000000000000000000000000000;	//		nop
memory[5] <= 32'b00000000000000000000000000000000;	//		nop
memory[6] <= 32'b00001000000000000000000000010010;	//		j	loop
memory[7] <= 32'b00000000000000000000000000000000;	//		nop
memory[8] <= 32'b00000000000000000000000000000000;	//		nop
memory[9] <= 32'b00000000000000000000000000000000;	//		nop
memory[10] <= 32'b00000000000000000000000000000000;	//		nop
memory[11] <= 32'b00000000000000000000000000000000;	//		nop
memory[12] <= 32'b00100000000010011111111111111111;	//		addi	$t1, $0, -1
memory[13] <= 32'b00000000000000000000000000000000;	//		nop
memory[14] <= 32'b00000000000000000000000000000000;	//		nop
memory[15] <= 32'b00000000000000000000000000000000;	//		nop
memory[16] <= 32'b00000000000000000000000000000000;	//		nop
memory[17] <= 32'b00000000000000000000000000000000;	//		nop
memory[18] <= 32'b00100001000010000000000000001010;	//	loop:	addi	$t0, $t0, 10
memory[19] <= 32'b00000000000000000000000000000000;	//		nop
memory[20] <= 32'b00000000000000000000000000000000;	//		nop
memory[21] <= 32'b00000000000000000000000000000000;	//		nop
memory[22] <= 32'b00000000000000000000000000000000;	//		nop
memory[23] <= 32'b00000000000000000000000000000000;	//		nop
memory[24] <= 32'b00001100000000000000000000101010;	//		jal	loop1
memory[25] <= 32'b00000000000000000000000000000000;	//		nop
memory[26] <= 32'b00000000000000000000000000000000;	//		nop
memory[27] <= 32'b00000000000000000000000000000000;	//		nop
memory[28] <= 32'b00000000000000000000000000000000;	//		nop
memory[29] <= 32'b00000000000000000000000000000000;	//		nop
memory[30] <= 32'b00100000000010000000000001100100;	//		addi	$t0, $0, 100
memory[31] <= 32'b00000000000000000000000000000000;	//		nop
memory[32] <= 32'b00000000000000000000000000000000;	//		nop
memory[33] <= 32'b00000000000000000000000000000000;	//		nop
memory[34] <= 32'b00000000000000000000000000000000;	//		nop
memory[35] <= 32'b00000000000000000000000000000000;	//		nop
memory[36] <= 32'b00001000000000000000000000110110;	//		j	exit
memory[37] <= 32'b00000000000000000000000000000000;	//		nop
memory[38] <= 32'b00000000000000000000000000000000;	//		nop
memory[39] <= 32'b00000000000000000000000000000000;	//		nop
memory[40] <= 32'b00000000000000000000000000000000;	//		nop
memory[41] <= 32'b00000000000000000000000000000000;	//		nop
memory[42] <= 32'b00100001000010000000000000001010;	//	loop1:	addi	$t0, $t0, 10
memory[43] <= 32'b00000000000000000000000000000000;	//		nop
memory[44] <= 32'b00000000000000000000000000000000;	//		nop
memory[45] <= 32'b00000000000000000000000000000000;	//		nop
memory[46] <= 32'b00000000000000000000000000000000;	//		nop
memory[47] <= 32'b00000000000000000000000000000000;	//		nop
memory[48] <= 32'b00000011111000000000000000001000;	//		jr	$ra
memory[49] <= 32'b00000000000000000000000000000000;	//		nop
memory[50] <= 32'b00000000000000000000000000000000;	//		nop
memory[51] <= 32'b00000000000000000000000000000000;	//		nop
memory[52] <= 32'b00000000000000000000000000000000;	//		nop
memory[53] <= 32'b00000000000000000000000000000000;	//		nop
memory[54] <= 32'b00100001000010000000000001100100;	//	exit:	addi	$t0, $t0, 100
memory[55] <= 32'b00000000000000000000000000000000;	//		nop
memory[56] <= 32'b00000000000000000000000000000000;	//		nop
memory[57] <= 32'b00000000000000000000000000000000;	//		nop
memory[58] <= 32'b00000000000000000000000000000000;	//		nop
memory[59] <= 32'b00000000000000000000000000000000;	//		nop
*/

/* //BRANCH TESTING
memory[0] <= 32'b00100000000010000000000000000001;	//			addi	$t0, $0, 1
memory[1] <= 32'b00000000000000000000000000000000;	//			nop
memory[2] <= 32'b00000000000000000000000000000000;	//			nop
memory[3] <= 32'b00000000000000000000000000000000;	//			nop
memory[4] <= 32'b00000000000000000000000000000000;	//			nop
memory[5] <= 32'b00000000000000000000000000000000;	//			nop
memory[6] <= 32'b00000101000000000000000000110101;	//			bltz	$t0, wrongBLTZ
memory[7] <= 32'b00000000000000000000000000000000;	//			nop
memory[8] <= 32'b00000000000000000000000000000000;	//			nop
memory[9] <= 32'b00000000000000000000000000000000;	//			nop
memory[10] <= 32'b00000000000000000000000000000000;	//			nop
memory[11] <= 32'b00000000000000000000000000000000;	//			nop
memory[12] <= 32'b00011001000000000000000000110101;	//			blez	$t0, wrongBLEZ
memory[13] <= 32'b00000000000000000000000000000000;	//			nop
memory[14] <= 32'b00000000000000000000000000000000;	//			nop
memory[15] <= 32'b00000000000000000000000000000000;	//			nop
memory[16] <= 32'b00000000000000000000000000000000;	//			nop
memory[17] <= 32'b00000000000000000000000000000000;	//			nop
memory[18] <= 32'b00100000000010011111111111111111;	//			addi	$t1, $0, -1
memory[19] <= 32'b00000000000000000000000000000000;	//			nop
memory[20] <= 32'b00000000000000000000000000000000;	//			nop
memory[21] <= 32'b00000000000000000000000000000000;	//			nop
memory[22] <= 32'b00000000000000000000000000000000;	//			nop
memory[23] <= 32'b00000000000000000000000000000000;	//			nop
memory[24] <= 32'b00011101001000000000000000101111;	//			bgtz	$t1, wrongBGTZ
memory[25] <= 32'b00000000000000000000000000000000;	//			nop
memory[26] <= 32'b00000000000000000000000000000000;	//			nop
memory[27] <= 32'b00000000000000000000000000000000;	//			nop
memory[28] <= 32'b00000000000000000000000000000000;	//			nop
memory[29] <= 32'b00000000000000000000000000000000;	//			nop
memory[30] <= 32'b00000101001000010000000000101111;	//			bgez	$t1, wrongBGEZ
memory[31] <= 32'b00000000000000000000000000000000;	//			nop
memory[32] <= 32'b00000000000000000000000000000000;	//			nop
memory[33] <= 32'b00000000000000000000000000000000;	//			nop
memory[34] <= 32'b00000000000000000000000000000000;	//			nop
memory[35] <= 32'b00000000000000000000000000000000;	//			nop
memory[36] <= 32'b00010001000010010000000000101111;	//			beq	$t0, $t1, wrongBEQ
memory[37] <= 32'b00000000000000000000000000000000;	//			nop
memory[38] <= 32'b00000000000000000000000000000000;	//			nop
memory[39] <= 32'b00000000000000000000000000000000;	//			nop
memory[40] <= 32'b00000000000000000000000000000000;	//			nop
memory[41] <= 32'b00000000000000000000000000000000;	//			nop
memory[42] <= 32'b00100000000010010000000000000001;	//			addi	$t1, $0, 1
memory[43] <= 32'b00000000000000000000000000000000;	//			nop
memory[44] <= 32'b00000000000000000000000000000000;	//			nop
memory[45] <= 32'b00000000000000000000000000000000;	//			nop
memory[46] <= 32'b00000000000000000000000000000000;	//			nop
memory[47] <= 32'b00000000000000000000000000000000;	//			nop
memory[48] <= 32'b00010101000010010000000000101001;	//			bne	$t0, $t1, wrongBNE
memory[49] <= 32'b00000000000000000000000000000000;	//			nop
memory[50] <= 32'b00000000000000000000000000000000;	//			nop
memory[51] <= 32'b00000000000000000000000000000000;	//			nop
memory[52] <= 32'b00000000000000000000000000000000;	//			nop
memory[53] <= 32'b00000000000000000000000000000000;	//			nop
memory[54] <= 32'b00010001000010010000000000101001;	//			beq	$t0, $t1, rightBEQ
memory[55] <= 32'b00000000000000000000000000000000;	//			nop
memory[56] <= 32'b00000000000000000000000000000000;	//			nop
memory[57] <= 32'b00000000000000000000000000000000;	//			nop
memory[58] <= 32'b00000000000000000000000000000000;	//			nop
memory[59] <= 32'b00000000000000000000000000000000;	//			nop
memory[60] <= 32'b00100000000010101111111111110110;	//	wrongBLTZ:	addi	$t2, $0, -10
memory[61] <= 32'b00000000000000000000000000000000;	//			nop
memory[62] <= 32'b00000000000000000000000000000000;	//			nop
memory[63] <= 32'b00000000000000000000000000000000;	//			nop
memory[64] <= 32'b00000000000000000000000000000000;	//			nop
memory[65] <= 32'b00000000000000000000000000000000;	//			nop
memory[66] <= 32'b00100000000010101111111111101100;	//	wrongBLEZ:	addi	$t2, $0, -20
memory[67] <= 32'b00000000000000000000000000000000;	//			nop
memory[68] <= 32'b00000000000000000000000000000000;	//			nop
memory[69] <= 32'b00000000000000000000000000000000;	//			nop
memory[70] <= 32'b00000000000000000000000000000000;	//			nop
memory[71] <= 32'b00000000000000000000000000000000;	//			nop
memory[72] <= 32'b00100000000010101111111111100010;	//	wrongBGTZ:	addi	$t2, $0, -30
memory[73] <= 32'b00000000000000000000000000000000;	//			nop
memory[74] <= 32'b00000000000000000000000000000000;	//			nop
memory[75] <= 32'b00000000000000000000000000000000;	//			nop
memory[76] <= 32'b00000000000000000000000000000000;	//			nop
memory[77] <= 32'b00000000000000000000000000000000;	//			nop
memory[78] <= 32'b00100000000010101111111111011000;	//	wrongBGEZ:	addi	$t2, $0, -40
memory[79] <= 32'b00000000000000000000000000000000;	//			nop
memory[80] <= 32'b00000000000000000000000000000000;	//			nop
memory[81] <= 32'b00000000000000000000000000000000;	//			nop
memory[82] <= 32'b00000000000000000000000000000000;	//			nop
memory[83] <= 32'b00000000000000000000000000000000;	//			nop
memory[84] <= 32'b00100000000010101111111111001110;	//	wrongBEQ:	addi	$t2, $0, -50
memory[85] <= 32'b00000000000000000000000000000000;	//			nop
memory[86] <= 32'b00000000000000000000000000000000;	//			nop
memory[87] <= 32'b00000000000000000000000000000000;	//			nop
memory[88] <= 32'b00000000000000000000000000000000;	//			nop
memory[89] <= 32'b00000000000000000000000000000000;	//			nop
memory[90] <= 32'b00100000000010101111111111000100;	//	wrongBNE:	addi	$t2, $0, -60
memory[91] <= 32'b00000000000000000000000000000000;	//			nop
memory[92] <= 32'b00000000000000000000000000000000;	//			nop
memory[93] <= 32'b00000000000000000000000000000000;	//			nop
memory[94] <= 32'b00000000000000000000000000000000;	//			nop
memory[95] <= 32'b00000000000000000000000000000000;	//			nop
memory[96] <= 32'b00100000000010000000000000000000;	//	rightBEQ:	addi	$t0, $0, 0
memory[97] <= 32'b00000000000000000000000000000000;	//			nop
memory[98] <= 32'b00000000000000000000000000000000;	//			nop
memory[99] <= 32'b00000000000000000000000000000000;	//			nop
memory[100] <= 32'b00000000000000000000000000000000;	//			nop
memory[101] <= 32'b00000000000000000000000000000000;	//			nop
memory[102] <= 32'b00010101000010010000000000001011;	//			bne	$t0, $t1, rightBNE
memory[103] <= 32'b00000000000000000000000000000000;	//			nop
memory[104] <= 32'b00000000000000000000000000000000;	//			nop
memory[105] <= 32'b00000000000000000000000000000000;	//			nop
memory[106] <= 32'b00000000000000000000000000000000;	//			nop
memory[107] <= 32'b00000000000000000000000000000000;	//			nop
memory[108] <= 32'b00100000000010101111111110111010;	//			addi	$t2, $0, -70
memory[109] <= 32'b00000000000000000000000000000000;	//			nop
memory[110] <= 32'b00000000000000000000000000000000;	//			nop
memory[111] <= 32'b00000000000000000000000000000000;	//			nop
memory[112] <= 32'b00000000000000000000000000000000;	//			nop
memory[113] <= 32'b00000000000000000000000000000000;	//			nop
memory[114] <= 32'b00000101000000010000000000001011;	//	rightBNE:	bgez	$t0, rightBGEZ
memory[115] <= 32'b00000000000000000000000000000000;	//			nop
memory[116] <= 32'b00000000000000000000000000000000;	//			nop
memory[117] <= 32'b00000000000000000000000000000000;	//			nop
memory[118] <= 32'b00000000000000000000000000000000;	//			nop
memory[119] <= 32'b00000000000000000000000000000000;	//			nop
memory[120] <= 32'b00100000000010101111111110110000;	//			addi	$t2, $0, -80
memory[121] <= 32'b00000000000000000000000000000000;	//			nop
memory[122] <= 32'b00000000000000000000000000000000;	//			nop
memory[123] <= 32'b00000000000000000000000000000000;	//			nop
memory[124] <= 32'b00000000000000000000000000000000;	//			nop
memory[125] <= 32'b00000000000000000000000000000000;	//			nop
memory[126] <= 32'b00011001000000000000000000001011;	//	rightBGEZ:	blez	$t0, rightBLEZ
memory[127] <= 32'b00000000000000000000000000000000;	//			nop
memory[128] <= 32'b00000000000000000000000000000000;	//			nop
memory[129] <= 32'b00000000000000000000000000000000;	//			nop
memory[130] <= 32'b00000000000000000000000000000000;	//			nop
memory[131] <= 32'b00000000000000000000000000000000;	//			nop
memory[132] <= 32'b00100000000010101111111110100110;	//			addi	$t2, $0, -90
memory[133] <= 32'b00000000000000000000000000000000;	//			nop
memory[134] <= 32'b00000000000000000000000000000000;	//			nop
memory[135] <= 32'b00000000000000000000000000000000;	//			nop
memory[136] <= 32'b00000000000000000000000000000000;	//			nop
memory[137] <= 32'b00000000000000000000000000000000;	//			nop
memory[138] <= 32'b00011101001000000000000000001011;	//	rightBLEZ:	bgtz	$t1, rightBGTZ
memory[139] <= 32'b00000000000000000000000000000000;	//			nop
memory[140] <= 32'b00000000000000000000000000000000;	//			nop
memory[141] <= 32'b00000000000000000000000000000000;	//			nop
memory[142] <= 32'b00000000000000000000000000000000;	//			nop
memory[143] <= 32'b00000000000000000000000000000000;	//			nop
memory[144] <= 32'b00100000000010101111111110011100;	//			addi	$t2, $0, -100
memory[145] <= 32'b00000000000000000000000000000000;	//			nop
memory[146] <= 32'b00000000000000000000000000000000;	//			nop
memory[147] <= 32'b00000000000000000000000000000000;	//			nop
memory[148] <= 32'b00000000000000000000000000000000;	//			nop
memory[149] <= 32'b00000000000000000000000000000000;	//			nop
memory[150] <= 32'b00100000000010011111111111111111;	//	rightBGTZ:	addi	$t1, $0, -1
memory[151] <= 32'b00000000000000000000000000000000;	//			nop
memory[152] <= 32'b00000000000000000000000000000000;	//			nop
memory[153] <= 32'b00000000000000000000000000000000;	//			nop
memory[154] <= 32'b00000000000000000000000000000000;	//			nop
memory[155] <= 32'b00000000000000000000000000000000;	//			nop
memory[156] <= 32'b00000101001000000000000000001011;	//			bltz	$t1, rightBLTZ
memory[157] <= 32'b00000000000000000000000000000000;	//			nop
memory[158] <= 32'b00000000000000000000000000000000;	//			nop
memory[159] <= 32'b00000000000000000000000000000000;	//			nop
memory[160] <= 32'b00000000000000000000000000000000;	//			nop
memory[161] <= 32'b00000000000000000000000000000000;	//			nop
memory[162] <= 32'b00100000000010101111111110010010;	//			addi	$t2, $0, -110
memory[163] <= 32'b00000000000000000000000000000000;	//			nop
memory[164] <= 32'b00000000000000000000000000000000;	//			nop
memory[165] <= 32'b00000000000000000000000000000000;	//			nop
memory[166] <= 32'b00000000000000000000000000000000;	//			nop
memory[167] <= 32'b00000000000000000000000000000000;	//			nop
memory[168] <= 32'b00100000000010000000000001100100;	//	rightBLTZ:	addi	$t0, $0, 100
memory[169] <= 32'b00000000000000000000000000000000;	//			nop
memory[170] <= 32'b00000000000000000000000000000000;	//			nop
memory[171] <= 32'b00000000000000000000000000000000;	//			nop
memory[172] <= 32'b00000000000000000000000000000000;	//			nop
memory[173] <= 32'b00000000000000000000000000000000;	//			nop
memory[174] <= 32'b00100000000010010000000001100100;	//			addi	$t1, $0, 100
memory[175] <= 32'b00000000000000000000000000000000;	//			nop
memory[176] <= 32'b00000000000000000000000000000000;	//			nop
memory[177] <= 32'b00000000000000000000000000000000;	//			nop
memory[178] <= 32'b00000000000000000000000000000000;	//			nop
memory[179] <= 32'b00000000000000000000000000000000;	//			nop
memory[180] <= 32'b00100000000010100000000001100100;	//			addi	$t2, $0, 100
*/ 

//tested data forwarding
//memory[1] <= 32'b00100000000100010000000000000001;	//		addi	$s1, $zero, 1
//memory[2] <= 32'b00100000000100100000000000000010;	//		addi	$s2, $zero, 2
//memory[3] <= 32'b00100000000100110000000000000011;	//		addi	$s3, $zero, 3
//memory[4] <= 32'b00100000000101000000000000000100;	//		addi	$s4, $zero, 4memory[4] <= 32'b00000000000000000000000000000000;	//		nop
//memory[5] <= 32'b00000000000000000000000000000000;	//		nop
//memory[6] <= 32'b00000000000000000000000000000000;	//		nop
//memory[7] <= 32'b00000000000000000000000000000000;	//		nop
//memory[8] <= 32'b00000010010100011001100000100010;	//		sub	$s3, $s2, $s1
//memory[9] <= 32'b00000010011100011010000000100100;	//		and	$s4, $s3, $s1
//memory[10] <= 32'b00000000000000000000000000000000;	//		nop
//memory[11] <= 32'b00000000000000000000000000000000;	//		nop
//memory[12] <= 32'b00000000000000000000000000000000;	//		nop
//memory[13] <= 32'b00000000000000000000000000000000;	//		nop
//memory[14] <= 32'b00000010010100011001100000100010;	//		sub	$s3, $s2, $s1
//memory[15] <= 32'b00000010001100111010000000100100;	//		and	$s4, $s1, $s3
//memory[16] <= 32'b00000000000000000000000000000000;	//		nop
//memory[17] <= 32'b00000000000000000000000000000000;	//		nop
//memory[18] <= 32'b00000000000000000000000000000000;	//		nop
//memory[19] <= 32'b00000000000000000000000000000000;	//		nop
//memory[20] <= 32'b00000010010100011001100000100010;	//		sub	$s3, $s2, $s1
//memory[21] <= 32'b00100000000101010000000000000100;	//		addi	$s5, $zero, 4
//memory[22] <= 32'b00000010011100011010000000100100;	//		and	$s4, $s3, $s1
//memory[23] <= 32'b00000000000000000000000000000000;	//		nop
//memory[24] <= 32'b00000000000000000000000000000000;	//		nop
//memory[25] <= 32'b00000000000000000000000000000000;	//		nop
//memory[26] <= 32'b00000000000000000000000000000000;	//		nop
//memory[27] <= 32'b00000010010100011001100000100010;	//		sub	$s3, $s2, $s1
//memory[28] <= 32'b00100000000101010000000000000100;	//		addi	$s5, $zero, 4
//memory[29] <= 32'b00000010001100111010000000100100;	//		and	$s4, $s1, $s3
//memory[30] <= 32'b00000000000000000000000000000000;	//		nop
//memory[31] <= 32'b00000000000000000000000000000000;	//		nop
//memory[32] <= 32'b00000000000000000000000000000000;	//		nop
//memory[33] <= 32'b00100000000100010000000000000001;	//		addi	$s1, $zero, 1
//memory[34] <= 32'b00100000000100100000000000000010;	//		addi	$s2, $zero, 2
//memory[35] <= 32'b00100000000100110000000000000011;	//		addi	$s3, $zero, 3
//memory[36] <= 32'b00100000000101000000000000000100;	//		addi	$s4, $zero, 4
//memory[37] <= 32'b00000000000000000000000000000000;	//		nop
//memory[38] <= 32'b00000000000000000000000000000000;	//		nop
//memory[39] <= 32'b00000000000000000000000000000000;	//		nop
//memory[40] <= 32'b00000000000000000000000000000000;	//		nop
//memory[41] <= 32'b00000010010100111000100000100000;	//		add	$s1, $s2, $s3
//memory[42] <= 32'b00000010010101001000100000100000;	//		add	$s1, $s2, $s4
//memory[43] <= 32'b00000010001101001001100000100000;	//		add	$s3, $s1, $s4
//memory[44] <= 32'b00000000000000000000000000000000;	//		nop
//memory[45] <= 32'b00000000000000000000000000000000;	//		nop
//memory[46] <= 32'b00000000000000000000000000000000;	//		nop
//memory[47] <= 32'b00000000000000000000000000000000;	//		nop
//memory[48] <= 32'b00100000000100010000000000000001;	//		addi	$s1, $zero, 1
//memory[49] <= 32'b00100000000100100000000000000010;	//		addi	$s2, $zero, 2
//memory[50] <= 32'b00100000000100110000000000000011;	//		addi	$s3, $zero, 3
//memory[51] <= 32'b00100000000101000000000000000100;	//		addi	$s4, $zero, 4
//memory[52] <= 32'b00000000000000000000000000000000;	//		nop
//memory[53] <= 32'b00000000000000000000000000000000;	//		nop
//memory[54] <= 32'b00000000000000000000000000000000;	//		nop
//memory[55] <= 32'b00000000000000000000000000000000;	//		nop
//memory[56] <= 32'b00000010010100111000100000100000;	//		add	$s1, $s2, $s3
//memory[57] <= 32'b00000010010100011001100000100000;	//		add	$s3, $s2, $s1
//memory[58] <= 32'b00000010001100011000100000100010;	//		sub	$s1, $s1, $s1
//memory[59] <= 32'b00000000000000000000000000000000;	//		nop
//memory[60] <= 32'b00000000000000000000000000000000;	//		nop
//memory[61] <= 32'b00000000000000000000000000000000;	//		nop
//memory[62] <= 32'b00000000000000000000000000000000;	//		nop
//memory[63] <= 32'b00100000000100010000000000000001;	//		addi	$s1, $zero, 1
//memory[64] <= 32'b00100000000100100000000000000010;	//		addi	$s2, $zero, 2
//memory[65] <= 32'b00100000000100110000000000000011;	//		addi	$s3, $zero, 3
//memory[66] <= 32'b00100000000101000000000000000100;	//		addi	$s4, $zero, 4
//memory[67] <= 32'b00000000000000000000000000000000;	//		nop
//memory[68] <= 32'b00000000000000000000000000000000;	//		nop
//memory[69] <= 32'b00000000000000000000000000000000;	//		nop
//memory[70] <= 32'b00000000000000000000000000000000;	//		nop
//memory[71] <= 32'b00000010010100111000100000100000;	//		add	$s1, $s2, $s3
//memory[72] <= 32'b00000010010100111010000000100000;	//		add	$s4, $s2, $s3
//memory[73] <= 32'b00000010010100111010000000100000;	//		add	$s4, $s2, $s3
//memory[74] <= 32'b00000010001100101010100000100000;	//	    add $s5, $s1, $s2


//1 to 4 dependency 
//memory[0] <= 32'b00100000000100010000000000000001;    //        addi    $s1, $zero, 1
//memory[1] <= 32'b00100000000100100000000000000010;    //        addi    $s2, $zero, 2
//memory[2] <= 32'b00100000000100110000000000000011;    //        addi    $s3, $zero, 3
//memory[3] <= 32'b00100000000101000000000000000100;    //        addi    $s4, $zero, 4
//memory[4] <= 32'b00100000000101010000000000000101;    //        addi    $s5, $zero, 5
//memory[5] <= 32'b00100000000101100000000000000110;    //        addi    $s6, $zero, 6
//memory[6] <= 32'b00000000000000000000000000000000;    //        nop
//memory[7] <= 32'b00000000000000000000000000000000;    //        nop
//memory[8] <= 32'b00000000000000000000000000000000;    //        nop
//memory[9] <= 32'b00000000000000000000000000000000;    //        nop
//memory[10] <= 32'b00000010010100111000100000100000;    //        add    $s1, $s2, $s3
//memory[11] <= 32'b00100000000100100000000000000010;    //        addi    $s2, $zero, 2
//memory[12] <= 32'b00100000000100110000000000000011;    //        addi    $s3, $zero, 3
//memory[13] <= 32'b00000010001100101010000000100000;    //        add    $s4, $s1, $s2

//RAW
//memory[0] <= 32'b00100000000100010000000000000001;	//		addi	$s1, $zero, 1
//memory[1] <= 32'b00100000000100100000000000000010;	//		addi	$s2, $zero, 2
//memory[2] <= 32'b00100000000100110000000000000011;	//		addi	$s3, $zero, 3
//memory[3] <= 32'b00100000000101000000000000000100;	//		addi	$s4, $zero, 4
//memory[4] <= 32'b00000000000000000000000000000000;	//		nop
//memory[5] <= 32'b00000000000000000000000000000000;	//		nop
//memory[6] <= 32'b00000000000000000000000000000000;	//		nop
//memory[7] <= 32'b00000000000000000000000000000000;	//		nop
//memory[8] <= 32'b10101110100100010000000000000000;	//		sw	$s1, 0($s4)
//memory[9] <= 32'b10001110100101010000000000000000;	//		lw	$s5, 0($s4)
//memory[10] <= 32'b00000010101101001011000000100000;	//		add	$s6, $s5, $s4
memory[0] <= 32'b00100000000100010000000000000001;    //        addi    $s1, $0, 1
memory[1] <= 32'b00100000000100100000000000000001;    //        addi    $s2, $0, 1
memory[2] <= 32'b00000000000000000000000000000000;    //        nop
memory[3] <= 32'b00000000000000000000000000000000;    //        nop
memory[4] <= 32'b00000000000000000000000000000000;    //        nop
memory[5] <= 32'b00000000000000000000000000000000;    //        nop
memory[6] <= 32'b00010010001100100000000000000101;    //        beq    $s1, $s2, jump
memory[7] <= 32'b00000010001000000000000000010001;    //        mthi    $s1
memory[8] <= 32'b00000000000000000000000000000000;    //        nop
memory[9] <= 32'b00000000000000000000000000000000;    //        nop
memory[10] <= 32'b00000000000000000000000000000000;    //        nop
memory[11] <= 32'b00000000000000000000000000000000;    //        nop
memory[12] <= 32'b00100010001100010000000000001010;    //    jump:    addi    $s1, $s1, 10
//memory[0] <= 32'b00100000000100010000000001100100;    //        addi    $s1, $0, 100
//memory[1] <= 32'b00000000000000000000000000000000;    //        nop
//memory[2] <= 32'b00000000000000000000000000000000;    //        nop
//memory[3] <= 32'b00000000000000000000000000000000;    //        nop
//memory[4] <= 32'b00000000000000000000000000000000;    //        nop
//memory[5] <= 32'b00110110001100011010101010101010;    //        ori    $s1, $s1, 43690
//memory[6] <= 32'b00000000000000000000000000000000;    //        nop
//memory[7] <= 32'b00000000000100011000101010000000;    //        sll    $s1, $s1, 10
//memory[8] <= 32'b00100000000001000000000000000000;    //        addi    $a0, $0, 0
//memory[9] <= 32'b00100000000100000000000000000010;    //        addi    $s0, $0, 2
//memory[10] <= 32'b10101100100100000000000000000100;    //        sw    $s0, 4($a0)
//memory[11] <= 32'b10001100100100000000000000000100;    //        lw    $s0, 4($a0)








//memory[0] <= 32'b00110100000100100000000000000000; // main: ori $s2, $zero, 0
//memory[1] <= 32'b10001110010100100000000000000000; // lw $s2, 0($s2)
//memory[2] <= 32'b00110100000100110000000000000000; // ori $s3, $zero, 0
//memory[3] <= 32'b10001110011100110000000000000100; // lw $s3, 4($s3)
//memory[4] <= 32'b00000010010100111000100000100000; // add $s1, $s2, $s3
//memory[5] <= 32'b00000010001100111010000000100010; // sub $s4, $s1, $s3
//memory[6] <= 32'b00000010001101001000100000100010; // sub $s1, $s1, $s4
//memory[7] <= 32'b01110010001100111010000000000010; // mul $s4, $s1, $s3
//memory[8] <= 32'b00000010001100111010000000100010; // sub $s4, $s1, $s3
//memory[9] <= 32'b00000010010100111000100000100000; // add $s1, $s2, $s3
//memory[10] <= 32'b01110010001101001011000000000010; // mul $s6, $s1, $s4
//memory[11] <= 32'b00000010100101101000100000100010; // sub $s1, $s4, $s6
//memory[12] <= 32'b00000010010101101000100000100000; // add $s1, $s2, $s6
//memory[13] <= 32'b00110110001100011010101010101010; // ori $s1, $s1, 43690
//memory[14] <= 32'b00000000000100011000101010000000; // sll $s1, $s1, 10
//memory[15] <= 32'b00100010001101010000000000000000; // addi $s5, $s1, 0
//memory[16] <= 32'b00100010101101110000000000000000; // addi $s7, $s5, 0

//memory[17] <= 32'b00110100000100100000000000011000; // ori $s2, $zero, 24

//memory[18] <= 32'b10001110010100010000000000000000; // lw $s1, 0($s2)

//memory[19] <= 32'b00000010001101011010000000100010; // sub $s4, $s1, $s5

//memory[20] <= 32'b00000010001101111011000000100100; // and $s6, $s1, $s7

//memory[21] <= 32'b00000010001101101011100000100101; // or $s7, $s1, $s6

//memory[22] <= 32'b00000010001100111001000000100010; // sub $s2, $s1, $s3

//memory[23] <= 32'b00000010010101010100000000100100; // and $t0, $s2, $s5

//memory[24] <= 32'b00000010110100100100100000100101; // or $t1, $s6, $s2

//memory[25] <= 32'b00000010010100100101000000100000; // add $t2, $s2, $s2

//memory[26] <= 32'b00110100000100010000000000000000; // ori $s1, $zero, 0

//memory[27] <= 32'b10101110001010010000000000000100; // sw $t1, 4($s1)

//memory[28] <= 32'b10001110001010100000000000000100; // lw $t2, 4($s1)

//memory[29] <= 32'b00000010001100111001000000100010; // sub $s2, $s1, $s3

//memory[30] <= 32'b00000010010101010101100000100101; // or $t3, $s2, $s5

//memory[31] <= 32'b00000010010100100110000000100000; // add $t4, $s2, $s2

//memory[32] <= 32'b00000010010100100101000000100101; // or $t2, $s2, $s2

//memory[33] <= 32'b00000010111010101010000000100000; // add $s4, $s7, $t2

//memory[34] <= 32'b00110100000010010000000000000000; // ori $t1, $zero, 0

//memory[35] <= 32'b10001101001010000000000000000000; // lw $t0, 0($t1)

//memory[36] <= 32'b10001101001010100000000000000100; // lw $t2, 4($t1)

//memory[37] <= 32'b10101101001010100000000000000000; // sw $t2, 0($t1)

//memory[38] <= 32'b10101101001010000000000000000100; // sw $t0, 4($t1)

//memory[39] <= 32'b10001101001010000000000000000000; // lw $t0, 0($t1)

//memory[40] <= 32'b10001101001010100000000000000100; // lw $t2, 4($t1)

//memory[41] <= 32'b00110100000001000000000000011000; // ori $a0, $zero, 24

//memory[42] <= 32'b00001000000000000000000000101101; // j start

//memory[43] <= 32'b00100000000001001111111111111111; // addi $a0, $zero, -1

//memory[44] <= 32'b00100000000001001111111111111111; // addi $a0, $zero, -1

//memory[45] <= 32'b10001100100100000000000000000100; // start: lw $s0, 4($a0)

//memory[46] <= 32'b10101100100100000000000000000000; // sw $s0, 0($a0)

//memory[47] <= 32'b00000110000000010000000000000011; // branch1: bgez $s0, branch2

//memory[48] <= 32'b00100010000100000000000000000001; // addi $s0, $s0, 1

//memory[49] <= 32'b00000110000000011111111111111101; // bgez $s0, branch1

//memory[50] <= 32'b00001000000000000000000000111101; // j error

//memory[51] <= 32'b00100000000100001111111111111111; // branch2: addi $s0, $zero, -1

//memory[52] <= 32'b00000110000000000000000000000011; // bltz $s0, branch3

//memory[53] <= 32'b00100000000100000000000000000001; // addi $s0, $zero, 1

//memory[54] <= 32'b00011110000000001111111111111100; // bgtz $s0, branch2

//memory[55] <= 32'b00001000000000000000000000111101; // j error

//memory[56] <= 32'b00000110000000000000000000000011; // branch3: bltz $s0, done

//memory[57] <= 32'b00100000000100001111111111111111; // addi $s0, $zero, -1

//memory[58] <= 32'b00000110000000001111111111111101; // bltz $s0, branch3

//memory[59] <= 32'b00001000000000000000000000111101; // j error

//memory[60] <= 32'b00001000000000000000000000111100; // done: j done

//memory[61] <= 32'b00001000000000000000000000111101; // error: j error  
    end
    
    always @ * begin
    Instruction = memory[Address[11:2]];
    end
    

endmodule